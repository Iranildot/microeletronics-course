* TASK 1 - INVERTER (MICROELETRONICS COURSE)

.SUBCKT inv IN OUT VDD GND
X0 OUT IN GND GND sky130_fd_pr__nfet_01v8 w=1000000u  l=150000u
X1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 w=3000000u l=150000u
.ENDS
