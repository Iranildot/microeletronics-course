magic
tech sky130A
timestamp 1730211546
<< metal4 >>
rect -2570 2300 0 2350
rect -2570 130 -170 2300
rect -50 130 0 2300
rect -2570 80 0 130
rect 80 2300 2650 2350
rect 80 130 2480 2300
rect 2600 130 2650 2300
rect 80 80 2650 130
rect -2570 -70 0 -20
rect -2570 -2240 -170 -70
rect -50 -2240 0 -70
rect -2570 -2290 0 -2240
rect 80 -70 2650 -20
rect 80 -2240 2480 -70
rect 2600 -2240 2650 -70
rect 80 -2290 2650 -2240
<< via4 >>
rect -170 130 -50 2300
rect 2480 130 2600 2300
rect -170 -2240 -50 -70
rect 2480 -2240 2600 -70
<< mimcap2 >>
rect -2550 2280 -320 2330
rect -2550 150 -2500 2280
rect -370 150 -320 2280
rect -2550 100 -320 150
rect 100 2280 2330 2330
rect 100 150 150 2280
rect 2280 150 2330 2280
rect 100 100 2330 150
rect -2550 -90 -320 -40
rect -2550 -2220 -2500 -90
rect -370 -2220 -320 -90
rect -2550 -2270 -320 -2220
rect 100 -90 2330 -40
rect 100 -2220 150 -90
rect 2280 -2220 2330 -90
rect 100 -2270 2330 -2220
<< mimcap2contact >>
rect -2500 150 -370 2280
rect 150 150 2280 2280
rect -2500 -2220 -370 -90
rect 150 -2220 2280 -90
<< metal5 >>
rect -190 2300 -30 2320
rect 2460 2300 2620 2320
rect -2520 2280 -350 2300
rect -2520 150 -2500 2280
rect -370 150 -350 2280
rect -2520 130 -350 150
rect -190 130 -170 2300
rect -50 130 -30 2300
rect 130 2280 2300 2300
rect 130 150 150 2280
rect 2280 150 2300 2280
rect 130 130 2300 150
rect 2460 130 2480 2300
rect 2600 130 2620 2300
rect -1565 -70 -1405 130
rect -190 -70 -30 130
rect 1085 -70 1245 130
rect 2460 -70 2620 130
rect -2520 -90 -350 -70
rect -2520 -2220 -2500 -90
rect -370 -2220 -350 -90
rect -2520 -2240 -350 -2220
rect -190 -2240 -170 -70
rect -50 -2240 -30 -70
rect 130 -90 2300 -70
rect 130 -2220 150 -90
rect 2280 -2220 2300 -90
rect 130 -2240 2300 -2220
rect 2460 -2240 2480 -70
rect 2600 -2240 2620 -70
rect -190 -2260 -30 -2240
rect 2460 -2260 2620 -2240
<< end >>
