* SPICE3 file created from lc_filter_pex_magic.ext - technology: sky130A

*.option scale=5000u

.subckt lc_filter_pex_magic p1 p2 gnd
X0 p1 p2 sky130_fd_pr__cap_mim_m3_2 l=22.3 w=22.3
X1 p1 p2 sky130_fd_pr__cap_mim_m3_2 l=22.3 w=22.3
X2 p1 p2 sky130_fd_pr__cap_mim_m3_2 l=22.3 w=22.3
X3 p1 p2 sky130_fd_pr__cap_mim_m3_2 l=22.3 w=22.3
C0 p1 p2 167.71fF
C1 p1 gnd 0.49fF
C2 p2 gnd 33.62fF
.ends
