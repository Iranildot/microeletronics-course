** sch_path: /home/isales/sky130_skel/xschem_sky130/MICRO/LC-LVS.sch

.subckt lc_filter_lvs_xschem p1 p2 gnd
XC1 p1 p2 sky130_fd_pr__cap_mim_m3_2 W=22.3 L=22.3 MF=4 m=4
R1 p1 p2 sky130_fd_pr__res_generic_m5 W=12 L=1 m=1
.ends
