* TASK 1 - INVERTER (MICROELETRONICS COURSE)

.option scale=1e-8

* INCLUDING SKY130 TECHNOLOGY
.lib "/edatools/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* INCLUDING THE INVERTER SUBCIRCUIT
.include ./INV_ideal.spice

* CREATING A 1.8 V DC POWER
Vdd VDD GND 1.8

* INSTANTIATING INVERTER
X1 IN OUT VDD GND inv

* CREATING A PULSE
Vin IN GND pulse(0 1.8 1p 10p 10p 1n 2n)

* PERFORMING SIMULATION AND PLOTTING
.tran 10e-12 2e-9

.control
run
plot IN OUT
.endc
.end

