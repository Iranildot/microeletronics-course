magic
tech sky130A
timestamp 1730212973
<< psubdiff >>
rect -11435 385 -10175 415
rect -11435 -815 -11405 385
rect -10205 -815 -10175 385
rect -11435 -845 -10175 -815
<< psubdiffcont >>
rect -11405 -815 -10205 385
<< locali >>
rect -11435 385 -10175 415
rect -11435 -815 -11405 385
rect -10205 -815 -10175 385
rect -11435 -845 -10175 -815
<< viali >>
rect -11405 -815 -10205 385
<< metal1 >>
rect -11435 385 -10175 415
rect -11435 -815 -11405 385
rect -10205 -815 -10175 385
rect -11435 -845 -10175 -815
<< via1 >>
rect -11405 -815 -10205 385
<< metal2 >>
rect -11435 385 -10175 415
rect -11435 -815 -11405 385
rect -10205 -815 -10175 385
rect -11435 -845 -10175 -815
<< via2 >>
rect -11405 -815 -10205 385
<< metal3 >>
rect -11435 385 -10175 415
rect -11435 -815 -11405 385
rect -10205 -815 -10175 385
rect -11435 -845 -10175 -815
<< metal4 >>
rect -7480 24 -7320 4560
rect -4830 24 -4670 4560
rect 6600 24 7800 1257
rect -7480 -1176 7800 24
rect -2360 -2375 -1160 -1176
<< metal5 >>
rect -2360 13200 -1160 14400
rect -7485 12000 1200 13200
rect -7485 9150 -7325 12000
rect -4835 9150 -4675 12000
use mim_cap_m4  mim_cap_m4_0
timestamp 1730211546
transform 1 0 -5917 0 1 6850
box -2570 -2290 2650 2350
use inductor  inductor_0
timestamp 1730208995
transform 1 0 -19600 0 1 -18400
box 19600 18400 31600 31600
<< end >>
