* SPICE3 file created from INV3.ext - technology: sky130A

.SUBCKT inv IN OUT VDD GND
M1000 OUT IN VDD w_n58_185# pshort_model.0 w=300 l=15
+  ad=11400 pd=676 as=11400 ps=676
M1001 OUT IN GND SUB nshort_model.0 w=100 l=15
+  ad=3800 pd=276 as=3800 ps=276
C0 IN GND 0.03fF
C1 OUT GND 0.08fF
C2 VDD GND 0.01fF
C3 OUT IN 0.04fF
C4 OUT w_n58_185# 0.00fF
C5 IN VDD 0.02fF
C6 OUT VDD 0.22fF
C7 w_n58_185# VDD 0.00fF
C8 GND SUB 0.39fF
C9 OUT SUB 0.10fF
C10 VDD SUB 0.39fF
C11 IN SUB 0.30fF
C12 w_n58_185# SUB 0.53fF
.ENDS
