magic
tech sky130A
timestamp 1729002766
<< nwell >>
rect -58 185 73 525
<< nmos >>
rect 0 20 15 120
<< pmos >>
rect 0 205 15 505
<< ndiff >>
rect -38 105 0 120
rect -38 80 -32 105
rect -15 80 0 105
rect -38 55 0 80
rect -38 30 -32 55
rect -15 30 0 55
rect -38 20 0 30
rect 15 110 53 120
rect 15 85 30 110
rect 47 85 53 110
rect 15 60 53 85
rect 15 35 30 60
rect 47 35 53 60
rect 15 20 53 35
<< pdiff >>
rect -38 492 0 505
rect -38 475 -32 492
rect -15 475 0 492
rect -38 457 0 475
rect -38 440 -32 457
rect -15 440 0 457
rect -38 422 0 440
rect -38 405 -32 422
rect -15 405 0 422
rect -38 387 0 405
rect -38 370 -32 387
rect -15 370 0 387
rect -38 352 0 370
rect -38 335 -32 352
rect -15 335 0 352
rect -38 317 0 335
rect -38 300 -32 317
rect -15 300 0 317
rect -38 282 0 300
rect -38 265 -32 282
rect -15 265 0 282
rect -38 247 0 265
rect -38 230 -32 247
rect -15 230 0 247
rect -38 205 0 230
rect 15 492 53 505
rect 15 475 30 492
rect 47 475 53 492
rect 15 457 53 475
rect 15 440 30 457
rect 47 440 53 457
rect 15 422 53 440
rect 15 405 30 422
rect 47 405 53 422
rect 15 387 53 405
rect 15 370 30 387
rect 47 370 53 387
rect 15 352 53 370
rect 15 335 30 352
rect 47 335 53 352
rect 15 317 53 335
rect 15 300 30 317
rect 47 300 53 317
rect 15 282 53 300
rect 15 265 30 282
rect 47 265 53 282
rect 15 247 53 265
rect 15 230 30 247
rect 47 230 53 247
rect 15 205 53 230
<< ndiffc >>
rect -32 80 -15 105
rect -32 30 -15 55
rect 30 85 47 110
rect 30 35 47 60
<< pdiffc >>
rect -32 475 -15 492
rect -32 440 -15 457
rect -32 405 -15 422
rect -32 370 -15 387
rect -32 335 -15 352
rect -32 300 -15 317
rect -32 265 -15 282
rect -32 230 -15 247
rect 30 475 47 492
rect 30 440 47 457
rect 30 405 47 422
rect 30 370 47 387
rect 30 335 47 352
rect 30 300 47 317
rect 30 265 47 282
rect 30 230 47 247
<< poly >>
rect 0 505 15 530
rect 0 175 15 205
rect -35 166 15 175
rect -35 149 -26 166
rect -9 149 15 166
rect -35 140 15 149
rect 0 120 15 140
rect 0 -5 15 20
<< polycont >>
rect -26 149 -9 166
<< locali >>
rect -43 560 -10 577
rect 7 560 25 577
rect 42 560 59 577
rect -32 492 -15 560
rect -32 457 -15 475
rect -32 422 -15 440
rect -32 387 -15 405
rect -32 352 -15 370
rect -32 317 -15 335
rect -32 282 -15 300
rect -32 247 -15 265
rect -32 210 -15 230
rect 30 492 47 500
rect 30 457 47 475
rect 30 422 47 440
rect 30 387 47 405
rect 30 352 47 370
rect 30 317 47 335
rect 30 282 47 300
rect 30 247 47 265
rect -35 166 0 175
rect -35 149 -26 166
rect -9 149 0 166
rect -35 140 0 149
rect -32 105 -15 115
rect -32 55 -15 80
rect -32 -35 -15 30
rect 30 110 47 230
rect 30 60 47 85
rect 30 25 47 35
rect -43 -52 -10 -35
rect 7 -52 24 -35
rect 41 -52 58 -35
<< viali >>
rect -60 560 -43 577
rect -10 560 7 577
rect 25 560 42 577
rect 59 560 76 577
rect -60 -52 -43 -35
rect -10 -52 7 -35
rect 24 -52 41 -35
rect 58 -52 75 -35
<< metal1 >>
rect -70 577 85 585
rect -70 560 -60 577
rect -43 560 -10 577
rect 7 560 25 577
rect 42 560 59 577
rect 76 560 85 577
rect -70 550 85 560
rect -70 -35 85 -25
rect -70 -52 -60 -35
rect -43 -52 -10 -35
rect 7 -52 24 -35
rect 41 -52 58 -35
rect 75 -52 85 -35
rect -70 -60 85 -52
<< end >>
